library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.imem.all;

package data is

   constant data : mem_block_t := (
      0 => (
         x"01", x"84", x"00", x"38", x"00", x"A0", x"00", x"50", x"00", x"04", 
         x"2A", x"FC", x"00", x"24", x"24", x"24", x"24", x"24", x"24", x"24", 
         x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", 
         x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", 
         x"24", x"24", x"EC", x"00", x"00", x"2C", x"00", x"00", x"00", x"08", 
         x"00", x"00", x"70", x"00", x"00", x"08", x"FF", x"50", x"00", x"00", 
         x"08", x"00", x"00", x"21", x"FF", x"10", x"00", x"00", x"08", x"00", 
         x"00", x"80", x"FF", x"00", x"21", x"00", x"08", x"00", x"00", x"21", 
         x"20", x"00", x"D0", x"00", x"08", x"00", x"00", x"70", x"00", x"00", 
         x"00", x"FF", x"00", x"03", x"F9", x"00", x"08", x"00", x"00", x"08", 
         x"00", x"00", x"08", x"00", x"FF", x"00", x"08", x"FF", x"FF", x"FF", 
         x"04", x"08", x"00", x"07", x"00", x"00", x"FF", x"00", x"01", x"FB", 
         x"01", x"08", x"00", x"06", x"00", x"03", x"FF", x"00", x"FD", x"01", 
         x"08", x"00", x"00", x"00", x"0A", x"00", x"21", x"01", x"21", x"00", 
         x"00", x"FC", x"01", x"08", x"FF", x"08", x"21", x"00", x"01", x"00", 
         x"FC", x"01", x"08", x"00", x"00", x"00", x"0D", x"FF", x"09", x"01", 
         x"A4", x"00", x"09", x"00", x"00", x"00", x"FB", x"01", x"08", x"00", 
         x"08", x"21", x"08", x"00", x"00", x"00", x"D0", x"FF", x"0A", x"13", 
         x"2D", x"11", x"00", x"0F", x"2D", x"C0", x"01", x"0B", x"00", x"09", 
         x"00", x"01", x"00", x"00", x"D0", x"FF", x"0A", x"F5", x"00", x"01", 
         x"00", x"D0", x"FF", x"0A", x"13", x"02", x"21", x"00", x"C0", x"40", 
         x"21", x"21", x"D0", x"FF", x"0A", x"F7", x"01", x"2D", x"03", x"00", 
         x"08", x"00", x"08", x"23", x"D9", x"21", x"30", x"00", x"62", x"01", 
         x"21", x"02", x"22", x"00", x"31", x"24", x"01", x"23", x"00", x"01", 
         x"FA", x"42", x"08", x"00", x"30", x"00", x"78", x"01", x"21", x"03", 
         x"1C", x"00", x"03", x"FC", x"FC", x"FF", x"02", x"0D", x"01", x"24", 
         x"06", x"FF", x"0A", x"30", x"F5", x"57", x"FC", x"FF", x"02", x"F5", 
         x"01", x"08", x"0A", x"10", x"00", x"40", x"26", x"42", x"26", x"40", 
         x"26", x"08", x"10", x"00", x"03", x"00", x"03", x"40", x"10", x"21", 
         x"01", x"2E", x"02", x"02", x"00", x"23", x"40", x"00", x"FF", x"43", 
         x"0B", x"03", x"03", x"F5", x"00", x"21", x"40", x"00", x"FF", x"43", 
         x"F7", x"03", x"08", x"00", x"05", x"00", x"04", x"21", x"08", x"00", 
         x"23", x"0D", x"00", x"2A", x"0C", x"23", x"21", x"21", x"01", x"00", 
         x"2A", x"FB", x"03", x"08", x"00", x"43", x"23", x"08", x"21", x"C4", 
         x"00", x"09", x"FF", x"C5", x"00", x"02", x"FF", x"C5", x"63", x"08", 
         x"C4", x"08", x"C4", x"14", x"08", x"15", x"FF", x"64", x"02", x"FF", 
         x"C4", x"25", x"02", x"00", x"C5", x"08", x"00", x"FF", x"E8", x"00", 
         x"02", x"FD", x"00", x"C4", x"08", x"C5", x"FF", x"C8", x"E8", x"00", 
         x"FF", x"FF", x"38", x"02", x"FA", x"00", x"20", x"E8", x"00", x"02", 
         x"FD", x"00", x"C5", x"00", x"03", x"FF", x"08", x"C4", x"08", x"C5", 
         x"C5", x"00", x"01", x"FF", x"25", x"03", x"C5", x"08", x"00", x"78", 
         x"00", x"C5", x"15", x"80", x"40", x"14", x"C4", x"21", x"80", x"21", 
         x"00", x"00", x"FF", x"21", x"25", x"01", x"FF", x"25", x"40", x"FF", 
         x"E8", x"21", x"FF", x"64", x"14", x"C4", x"00", x"04", x"00", x"90", 
         x"00", x"C4", x"14", x"00", x"08", x"18", x"E8", x"14", x"10", x"00", 
         x"00", x"08", x"01", x"FF", x"9B", x"01", x"FF", x"00", x"FB", x"FF", 
         x"14", x"10", x"08", x"18", x"D8", x"14", x"24", x"20", x"1C", x"18", 
         x"10", x"00", x"00", x"38", x"21", x"00", x"00", x"21", x"50", x"00", 
         x"EE", x"F4", x"61", x"0A", x"5B", x"08", x"55", x"00", x"9B", x"FF", 
         x"01", x"00", x"25", x"01", x"0D", x"4A", x"0E", x"F0", x"09", x"24", 
         x"38", x"25", x"11", x"25", x"23", x"EE", x"00", x"01", x"00", x"DD", 
         x"FF", x"57", x"E9", x"01", x"80", x"21", x"00", x"00", x"08", x"00", 
         x"11", x"5C", x"DD", x"00", x"9B", x"5C", x"01", x"00", x"DD", x"01", 
         x"24", x"20", x"1C", x"18", x"14", x"10", x"08", x"28", x"01", x"63", 
         x"76", x"01", x"64", x"2A", x"00", x"73", x"68", x"78", x"C5", x"00", 
         x"21", x"F4", x"A0", x"BE", x"21", x"EA", x"00", x"01", x"00", x"DC", 
         x"FF", x"56", x"B7", x"01", x"80", x"21", x"00", x"00", x"08", x"00", 
         x"EA", x"C4", x"53", x"00", x"EA", x"00", x"90", x"00", x"EA", x"C4", 
         x"C4", x"FC", x"04", x"24", x"EA", x"C4", x"44", x"62", x"9D", x"00", 
         x"21", x"E2", x"A0", x"BE", x"21", x"EA", x"00", x"9B", x"24", x"EA", 
         x"00", x"01", x"EA", x"14", x"03", x"EA", x"14", x"02", x"EA", x"14", 
         x"EA", x"14", x"05", x"EA", x"14", x"04", x"EA", x"14", x"07", x"EA", 
         x"14", x"06", x"EA", x"14", x"9B", x"23", x"EA", x"00", x"01", x"EA", 
         x"15", x"03", x"EA", x"15", x"02", x"EA", x"15", x"EA", x"15", x"05", 
         x"EA", x"15", x"04", x"EA", x"15", x"07", x"EA", x"15", x"06", x"EA", 
         x"15", x"BE", x"21", x"EA", x"00", x"9B", x"25", x"EA", x"00", x"9B", 
         x"FF", x"EA", x"00", x"FF", x"00", x"C8", x"02", x"C8", x"08", x"C9", 
         x"D0", x"28", x"00", x"24", x"20", x"1C", x"18", x"2C", x"14", x"21", 
         x"C4", x"FF", x"0D", x"08", x"00", x"80", x"FF", x"02", x"21", x"C8", 
         x"1F", x"C9", x"1D", x"00", x"27", x"00", x"F3", x"00", x"53", x"00", 
         x"C5", x"C4", x"80", x"40", x"21", x"80", x"21", x"21", x"40", x"21", 
         x"21", x"00", x"00", x"00", x"FF", x"FF", x"02", x"80", x"21", x"C8", 
         x"E3", x"C9", x"21", x"00", x"2C", x"21", x"24", x"28", x"20", x"1C", 
         x"18", x"14", x"08", x"30", x"9B", x"00", x"21", x"00", x"AC", x"01", 
         x"E0", x"14", x"FF", x"18", x"1C", x"10", x"09", x"FF", x"21", x"21", 
         x"9B", x"01", x"FF", x"2B", x"FB", x"21", x"1C", x"18", x"14", x"10", 
         x"08", x"20", x"C0", x"28", x"20", x"3C", x"38", x"34", x"30", x"2C", 
         x"24", x"1C", x"01", x"02", x"01", x"21", x"02", x"04", x"03", x"21", 
         x"21", x"00", x"FF", x"40", x"23", x"21", x"01", x"FD", x"FF", x"21", 
         x"27", x"FC", x"9B", x"10", x"00", x"BE", x"01", x"10", x"20", x"23", 
         x"E4", x"FF", x"04", x"FF", x"2B", x"2A", x"00", x"21", x"FF", x"64", 
         x"21", x"02", x"80", x"21", x"00", x"00", x"00", x"84", x"00", x"03", 
         x"00", x"E2", x"20", x"04", x"05", x"61", x"10", x"9B", x"DD", x"00", 
         x"BE", x"01", x"10", x"20", x"23", x"E4", x"FF", x"9B", x"DE", x"04", 
         x"05", x"61", x"FF", x"04", x"00", x"2B", x"D9", x"21", x"3C", x"38", 
         x"34", x"30", x"2C", x"28", x"24", x"20", x"1C", x"08", x"40", x"E0", 
         x"10", x"FF", x"FF", x"1C", x"18", x"14", x"FF", x"9B", x"FF", x"FE", 
         x"21", x"E4", x"FF", x"21", x"1C", x"18", x"14", x"10", x"9B", x"20", 
         x"D8", x"24", x"20", x"10", x"1C", x"21", x"18", x"14", x"03", x"01", 
         x"05", x"04", x"00", x"02", x"61", x"21", x"00", x"01", x"64", x"FF", 
         x"02", x"BB", x"C9", x"5B", x"CD", x"01", x"00", x"01", x"64", x"FF", 
         x"02", x"BA", x"BA", x"5B", x"20", x"00", x"01", x"02", x"01", x"FF", 
         x"64", x"FF", x"08", x"BE", x"FF", x"01", x"00", x"02", x"64", x"FF", 
         x"02", x"CC", x"CD", x"5B", x"B9", x"01", x"00", x"03", x"FF", x"2B", 
         x"12", x"21", x"FF", x"FF", x"00", x"64", x"21", x"9B", x"BA", x"21", 
         x"21", x"64", x"01", x"FF", x"9B", x"BA", x"2B", x"F2", x"00", x"00", 
         x"64", x"21", x"02", x"CD", x"BC", x"5B", x"C8", x"2B", x"21", x"24", 
         x"20", x"1C", x"18", x"14", x"10", x"07", x"21", x"61", x"28", x"E0", 
         x"14", x"21", x"04", x"1C", x"84", x"18", x"04", x"6F", x"FF", x"64", 
         x"23", x"00", x"14", x"C2", x"02", x"21", x"43", x"10", x"1C", x"18", 
         x"14", x"21", x"20", x"70", x"14", x"E0", x"18", x"21", x"04", x"14", 
         x"1C", x"84", x"21", x"01", x"01", x"00", x"02", x"21", x"21", x"02", 
         x"01", x"03", x"23", x"FF", x"FF", x"64", x"23", x"9B", x"20", x"04", 
         x"BE", x"00", x"FD", x"1C", x"18", x"14", x"20", x"FF", x"E4", x"20", 
         x"E8", x"14", x"10", x"21", x"02", x"01", x"00", x"01", x"21", x"21", 
         x"02", x"03", x"FF", x"64", x"FF", x"07", x"E4", x"FE", x"04", x"40", 
         x"23", x"14", x"10", x"20", x"FF", x"E4", x"18", x"D8", x"18", x"24", 
         x"20", x"1C", x"14", x"0C", x"00", x"22", x"21", x"21", x"01", x"41", 
         x"02", x"ED", x"00", x"0C", x"01", x"FF", x"2B", x"16", x"00", x"04", 
         x"80", x"21", x"00", x"21", x"00", x"00", x"14", x"21", x"EE", x"00", 
         x"EF", x"00", x"10", x"21", x"01", x"0C", x"FF", x"2B", x"ED", x"04", 
         x"24", x"20", x"1C", x"18", x"14", x"08", x"28", x"FA", x"01", x"0C", 
         x"3E", x"FF", x"04", x"03", x"FF", x"03", x"01", x"FA", x"03", x"FA", 
         x"03", x"03", x"00", x"03", x"FF", x"FA", x"03", x"04", x"00", x"FF", 
         x"FA", x"03", x"E8", x"14", x"56", x"00", x"02", x"0A", x"10", x"05", 
         x"68", x"14", x"00", x"08", x"18", x"14", x"D3", x"18", x"14", x"70", 
         x"D3", x"18", x"D8", x"20", x"00", x"24", x"10", x"1C", x"18", x"6F", 
         x"14", x"70", x"7C", x"7C", x"ED", x"50", x"7C", x"40", x"44", x"10", 
         x"04", x"68", x"FF", x"00", x"FF", x"FB", x"21", x"00", x"01", x"2B", 
         x"23", x"7C", x"ED", x"58", x"42", x"7C", x"40", x"44", x"10", x"01", 
         x"21", x"B5", x"7C", x"1F", x"00", x"4E", x"40", x"42", x"21", x"40", 
         x"10", x"44", x"56", x"01", x"20", x"F3", x"2B", x"24", x"20", x"1C", 
         x"18", x"14", x"10", x"60", x"D3", x"28", x"24", x"20", x"1C", x"18", 
         x"14", x"10", x"78", x"D3", x"28", x"18", x"21", x"04", x"06", x"21", 
         x"FF", x"3E", x"01", x"76", x"F8", x"F9", x"06", x"48", x"ED", x"7C", 
         x"02", x"6C", x"44", x"02", x"6C", x"FF", x"02", x"6C", x"FF", x"6C", 
         x"FF", x"1C", x"82", x"21", x"21", x"F7", x"7C", x"76", x"01", x"14", 
         x"00", x"68", x"00", x"21", x"3E", x"04", x"F6", x"21", x"44", x"00", 
         x"01", x"40", x"21", x"01", x"10", x"44", x"76", x"00", x"EE", x"00", 
         x"24", x"20", x"1C", x"18", x"14", x"10", x"00", x"28", x"D0", x"10", 
         x"00", x"2C", x"24", x"20", x"21", x"1C", x"21", x"28", x"18", x"6F", 
         x"14", x"70", x"64", x"82", x"64", x"40", x"10", x"44", x"1A", x"82", 
         x"00", x"21", x"00", x"21", x"31", x"7C", x"01", x"11", x"04", x"46", 
         x"21", x"00", x"F9", x"21", x"44", x"00", x"01", x"40", x"21", x"01", 
         x"44", x"10", x"04", x"F1", x"00", x"2C", x"28", x"24", x"20", x"1C", 
         x"18", x"14", x"10", x"08", x"30", x"C8", x"18", x"4D", x"2B", x"30", 
         x"34", x"2C", x"28", x"24", x"20", x"1C", x"14", x"10", x"51", x"21", 
         x"00", x"00", x"21", x"21", x"21", x"C0", x"06", x"00", x"6F", x"B4", 
         x"46", x"00", x"21", x"D0", x"21", x"4C", x"01", x"FF", x"01", x"16", 
         x"00", x"F4", x"21", x"04", x"06", x"64", x"FF", x"80", x"21", x"D0", 
         x"21", x"46", x"21", x"01", x"21", x"21", x"01", x"D0", x"FF", x"ED", 
         x"01", x"00", x"80", x"21", x"00", x"00", x"4D", x"21", x"21", x"C0", 
         x"06", x"98", x"B4", x"00", x"D0", x"00", x"25", x"01", x"FF", x"FF", 
         x"13", x"04", x"F6", x"21", x"14", x"06", x"64", x"FF", x"21", x"D0", 
         x"21", x"00", x"01", x"21", x"FF", x"D0", x"FF", x"01", x"EF", x"04", 
         x"34", x"30", x"2C", x"28", x"24", x"20", x"1C", x"18", x"14", x"10", 
         x"08", x"38", x"6C", x"21", x"95", x"21", x"D8", x"24", x"20", x"1C", 
         x"18", x"6F", x"14", x"00", x"70", x"50", x"00", x"70", x"3C", x"4B", 
         x"21", x"21", x"F0", x"F2", x"1B", x"97", x"00", x"01", x"00", x"0D", 
         x"00", x"13", x"00", x"F7", x"00", x"00", x"00", x"97", x"00", x"01", 
         x"00", x"F5", x"00", x"4D", x"02", x"00", x"B3", x"4B", x"21", x"CD", 
         x"00", x"4D", x"4B", x"21", x"CD", x"00", x"D8", x"24", x"20", x"1C", 
         x"18", x"14", x"6F", x"10", x"56", x"00", x"00", x"03", x"10", x"30", 
         x"12", x"00", x"D3", x"80", x"39", x"00", x"24", x"21", x"20", x"1C", 
         x"18", x"14", x"10", x"08", x"28", x"D3", x"88", x"00", x"00", x"70", 
         x"28", x"F0", x"F2", x"28", x"0D", x"01", x"97", x"00", x"01", x"00", 
         x"13", x"21", x"0D", x"00", x"F7", x"00", x"1B", x"00", x"1A", x"00", 
         x"0D", x"02", x"8A", x"00", x"14", x"00", x"62", x"18", x"14", x"00", 
         x"6B", x"18", x"14", x"00", x"E3", x"00", x"46", x"21", x"21", x"12", 
         x"01", x"30", x"00", x"14", x"00", x"BA", x"00", x"C0", x"A8", x"A8", 
         x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", 
         x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", 
         x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", 
         x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", 
         x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", 
         x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", 
         x"D0", x"DC", x"A8", x"A8", x"A8", x"E8", x"A8", x"A8", x"A8", x"F4", 
         x"A8", x"FC", x"A8", x"A8", x"A8", x"A8", x"08", x"A8", x"A8", x"A8", 
         x"A8", x"14", x"A8", x"20", x"54", x"A8", x"A8", x"A8", x"A8", x"A8", 
         x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", 
         x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", 
         x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", 
         x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", 
         x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", 
         x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"64", x"70", x"A8", x"A8", 
         x"A8", x"7C", x"A8", x"A8", x"A8", x"88", x"A8", x"90", x"A8", x"A8", 
         x"A8", x"A8", x"9C", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"B4", 
         x"41", x"52", x"00", x"78", x"20", x"00", x"00", x"64", x"6F", x"61", 
         x"20", x"32", x"00", x"72", x"2E", x"00", x"77", x"6D", x"20", x"74", 
         x"73", x"2E", x"00", x"6F", x"69", x"65", x"2E", x"00", x"20", x"6F", 
         x"00", x"73", x"65", x"79", x"00", x"20", x"64", x"00", x"64", x"20", 
         x"20", x"00", x"67", x"70", x"64", x"00", x"6F", x"6E", x"61", x"2E", 
         x"00", x"74", x"20", x"20", x"6F", x"6E", x"72", x"6D", x"69", x"2E", 
         x"00", x"73", x"20", x"73", x"6F", x"6E", x"2E", x"00", x"6C", x"6F", 
         x"72", x"20", x"73", x"6C", x"2E", x"00", x"6C", x"6F", x"72", x"20", 
         x"66", x"68", x"00", x"73", x"6C", x"20", x"6C", x"65", x"00", x"67", 
         x"69", x"65", x"65", x"61", x"6C", x"65", x"61", x"6D", x"72", x"00", 
         x"73", x"73", x"20", x"65", x"72", x"20", x"74", x"50", x"73", x"65", 
         x"72", x"00", x"73", x"73", x"74", x"61", x"20", x"68", x"68", x"20", 
         x"75", x"62", x"00", x"A1", x"00", x"00", x"00", x"B8", x"B4", x"B0", 
         x"DC", x"E8", x"04", x"00", x"40", x"00", x"00", x"00", x"60", x"00", 
         x"74", x"00", x"9C", x"00", x"B8", x"00", x"D8", x"00", x"F4", x"00", 
         x"0C", x"00", x"38", x"00", x"68", x"05", x"00", x"A8", x"00", x"00", 
         x"07", x"00", x"C4", x"00", x"9C", x"0F", x"00", x"18", x"00", x"00", 
         x"0F", x"00", x"24", x"00", x"00", x"06", x"00", x"34", x"00", x"BC", 
         x"C4", x"06", x"00", x"50", x"00", x"D4", x"C4", others => x"00"
      ),
      1 => (
         x"00", x"9D", x"00", x"3F", x"00", x"1E", x"00", x"1F", x"00", x"00", 
         x"08", x"FF", x"00", x"08", x"10", x"18", x"20", x"28", x"30", x"38", 
         x"40", x"48", x"50", x"58", x"60", x"68", x"70", x"78", x"80", x"88", 
         x"90", x"98", x"A0", x"A8", x"B0", x"B8", x"C0", x"C8", x"D0", x"D8", 
         x"F0", x"F8", x"05", x"00", x"00", x"00", x"00", x"00", x"20", x"00", 
         x"00", x"10", x"00", x"00", x"00", x"00", x"00", x"00", x"10", x"00", 
         x"00", x"00", x"10", x"10", x"00", x"00", x"00", x"00", x"00", x"00", 
         x"10", x"20", x"FF", x"00", x"10", x"00", x"00", x"00", x"10", x"10", 
         x"00", x"00", x"FF", x"00", x"00", x"00", x"10", x"00", x"00", x"00", 
         x"00", x"00", x"26", x"26", x"FF", x"00", x"00", x"00", x"F0", x"00", 
         x"00", x"F0", x"00", x"00", x"FF", x"40", x"00", x"00", x"00", x"FF", 
         x"40", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"FF", 
         x"00", x"00", x"00", x"00", x"2E", x"2E", x"FF", x"00", x"FF", x"00", 
         x"00", x"00", x"00", x"00", x"00", x"00", x"10", x"00", x"18", x"00", 
         x"00", x"FF", x"00", x"00", x"FF", x"00", x"10", x"00", x"00", x"00", 
         x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
         x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", 
         x"00", x"10", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", 
         x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
         x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"FF", x"00", x"00", 
         x"00", x"FF", x"00", x"00", x"00", x"00", x"10", x"00", x"38", x"10", 
         x"10", x"10", x"FF", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", 
         x"00", x"00", x"00", x"10", x"00", x"10", x"00", x"00", x"00", x"00", 
         x"10", x"00", x"00", x"80", x"00", x"28", x"00", x"28", x"00", x"00", 
         x"FF", x"30", x"00", x"00", x"00", x"00", x"00", x"00", x"10", x"00", 
         x"00", x"F0", x"01", x"FF", x"FF", x"FF", x"31", x"00", x"00", x"28", 
         x"28", x"00", x"00", x"00", x"FF", x"00", x"FF", x"FF", x"31", x"FF", 
         x"00", x"00", x"00", x"80", x"00", x"1B", x"10", x"1C", x"10", x"19", 
         x"10", x"00", x"80", x"24", x"24", x"2C", x"2C", x"20", x"00", x"10", 
         x"00", x"01", x"00", x"00", x"00", x"10", x"28", x"2C", x"FF", x"20", 
         x"00", x"2C", x"00", x"FF", x"00", x"10", x"28", x"2C", x"FF", x"20", 
         x"FF", x"2C", x"00", x"00", x"00", x"00", x"00", x"10", x"00", x"00", 
         x"28", x"00", x"00", x"10", x"00", x"30", x"10", x"20", x"00", x"14", 
         x"18", x"FF", x"14", x"00", x"00", x"01", x"20", x"00", x"10", x"81", 
         x"00", x"00", x"FF", x"81", x"00", x"00", x"FF", x"81", x"00", x"00", 
         x"81", x"00", x"81", x"80", x"00", x"80", x"00", x"00", x"00", x"00", 
         x"81", x"00", x"00", x"00", x"81", x"00", x"00", x"FF", x"1C", x"00", 
         x"00", x"FF", x"00", x"81", x"00", x"81", x"FF", x"00", x"1C", x"00", 
         x"FF", x"FF", x"FF", x"00", x"FF", x"00", x"1C", x"1C", x"00", x"00", 
         x"FF", x"00", x"81", x"00", x"00", x"FF", x"00", x"81", x"00", x"81", 
         x"81", x"00", x"00", x"00", x"00", x"00", x"81", x"00", x"00", x"01", 
         x"00", x"81", x"80", x"41", x"39", x"80", x"81", x"38", x"10", x"10", 
         x"32", x"2B", x"00", x"10", x"28", x"00", x"00", x"28", x"10", x"FF", 
         x"FF", x"10", x"FF", x"00", x"00", x"81", x"00", x"00", x"00", x"01", 
         x"00", x"81", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", 
         x"00", x"00", x"00", x"00", x"01", x"00", x"FF", x"00", x"FF", x"00", 
         x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", 
         x"00", x"00", x"00", x"00", x"88", x"00", x"00", x"80", x"1A", x"00", 
         x"01", x"18", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"00", 
         x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", 
         x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"FF", 
         x"00", x"00", x"FF", x"00", x"10", x"10", x"00", x"00", x"00", x"00", 
         x"00", x"00", x"FF", x"00", x"01", x"00", x"00", x"00", x"FF", x"00", 
         x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
         x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", 
         x"20", x"00", x"1E", x"01", x"20", x"01", x"00", x"00", x"00", x"FF", 
         x"00", x"00", x"FF", x"00", x"10", x"10", x"00", x"00", x"00", x"00", 
         x"01", x"81", x"01", x"00", x"01", x"00", x"01", x"00", x"01", x"81", 
         x"81", x"FF", x"00", x"10", x"01", x"81", x"00", x"00", x"FF", x"00", 
         x"20", x"00", x"1E", x"01", x"20", x"01", x"00", x"01", x"00", x"01", 
         x"00", x"00", x"01", x"80", x"00", x"01", x"80", x"00", x"01", x"80", 
         x"01", x"80", x"00", x"01", x"80", x"00", x"01", x"80", x"00", x"01", 
         x"80", x"00", x"01", x"80", x"01", x"00", x"01", x"00", x"00", x"01", 
         x"80", x"00", x"01", x"80", x"00", x"01", x"80", x"01", x"80", x"00", 
         x"01", x"80", x"00", x"01", x"80", x"00", x"01", x"80", x"00", x"01", 
         x"80", x"01", x"20", x"01", x"00", x"01", x"00", x"01", x"00", x"01", 
         x"00", x"01", x"00", x"FF", x"30", x"81", x"21", x"81", x"00", x"81", 
         x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"88", 
         x"1E", x"FF", x"00", x"00", x"30", x"00", x"00", x"11", x"20", x"81", 
         x"00", x"81", x"00", x"00", x"00", x"00", x"FF", x"00", x"01", x"00", 
         x"81", x"81", x"29", x"21", x"20", x"10", x"10", x"10", x"10", x"18", 
         x"10", x"00", x"00", x"30", x"FF", x"00", x"11", x"00", x"20", x"81", 
         x"FF", x"81", x"88", x"00", x"00", x"10", x"00", x"00", x"00", x"00", 
         x"00", x"00", x"00", x"00", x"01", x"00", x"10", x"00", x"02", x"00", 
         x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"80", x"20", 
         x"01", x"00", x"00", x"10", x"FF", x"20", x"00", x"00", x"00", x"00", 
         x"00", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
         x"00", x"00", x"00", x"00", x"00", x"A0", x"00", x"00", x"00", x"98", 
         x"88", x"00", x"00", x"00", x"B8", x"A8", x"00", x"FF", x"00", x"80", 
         x"03", x"FF", x"01", x"00", x"00", x"01", x"00", x"00", x"00", x"10", 
         x"02", x"00", x"00", x"00", x"10", x"00", x"00", x"28", x"00", x"01", 
         x"20", x"00", x"10", x"10", x"00", x"00", x"00", x"00", x"00", x"00", 
         x"00", x"FF", x"00", x"00", x"00", x"01", x"00", x"01", x"00", x"00", 
         x"01", x"00", x"00", x"00", x"10", x"02", x"00", x"01", x"00", x"00", 
         x"00", x"01", x"00", x"00", x"00", x"10", x"FF", x"28", x"00", x"00", 
         x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", 
         x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"01", x"00", x"FF", 
         x"20", x"02", x"00", x"20", x"00", x"00", x"00", x"00", x"01", x"00", 
         x"FF", x"00", x"00", x"00", x"00", x"80", x"00", x"00", x"00", x"00", 
         x"00", x"00", x"00", x"00", x"01", x"88", x"00", x"00", x"01", x"FF", 
         x"00", x"00", x"00", x"03", x"00", x"00", x"00", x"00", x"01", x"00", 
         x"00", x"00", x"00", x"03", x"00", x"00", x"00", x"00", x"00", x"00", 
         x"01", x"00", x"00", x"01", x"00", x"00", x"00", x"00", x"01", x"00", 
         x"00", x"00", x"00", x"03", x"00", x"00", x"00", x"00", x"00", x"10", 
         x"00", x"90", x"FF", x"00", x"00", x"01", x"28", x"01", x"00", x"28", 
         x"20", x"01", x"00", x"00", x"01", x"00", x"10", x"FF", x"00", x"00", 
         x"01", x"28", x"00", x"00", x"00", x"03", x"00", x"04", x"20", x"00", 
         x"00", x"00", x"00", x"00", x"00", x"00", x"28", x"01", x"00", x"FF", 
         x"00", x"80", x"00", x"00", x"00", x"00", x"00", x"01", x"00", x"00", 
         x"28", x"00", x"1E", x"27", x"00", x"28", x"28", x"00", x"00", x"00", 
         x"00", x"20", x"00", x"03", x"1E", x"FF", x"00", x"88", x"00", x"00", 
         x"00", x"00", x"80", x"00", x"00", x"00", x"00", x"20", x"28", x"00", 
         x"00", x"00", x"88", x"00", x"00", x"01", x"88", x"01", x"00", x"00", 
         x"01", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"02", x"00", 
         x"FF", x"00", x"00", x"80", x"00", x"00", x"00", x"00", x"20", x"28", 
         x"00", x"00", x"00", x"01", x"00", x"00", x"02", x"00", x"00", x"00", 
         x"28", x"00", x"00", x"00", x"00", x"02", x"00", x"FF", x"00", x"00", 
         x"00", x"00", x"00", x"00", x"00", x"00", x"88", x"80", x"00", x"04", 
         x"00", x"03", x"00", x"00", x"00", x"00", x"10", x"00", x"00", x"00", 
         x"10", x"10", x"00", x"20", x"00", x"00", x"00", x"28", x"FF", x"00", 
         x"FF", x"00", x"04", x"20", x"00", x"00", x"00", x"10", x"FF", x"00", 
         x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"02", x"00", x"00", 
         x"04", x"00", x"00", x"00", x"FF", x"00", x"00", x"02", x"00", x"02", 
         x"00", x"00", x"00", x"00", x"FF", x"02", x"00", x"00", x"00", x"FF", 
         x"02", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
         x"80", x"00", x"00", x"00", x"00", x"00", x"03", x"00", x"00", x"80", 
         x"03", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"01", 
         x"00", x"03", x"1E", x"1E", x"03", x"80", x"1E", x"80", x"80", x"04", 
         x"00", x"00", x"FF", x"8A", x"00", x"FF", x"88", x"01", x"00", x"10", 
         x"00", x"1E", x"03", x"80", x"9C", x"1E", x"80", x"80", x"04", x"00", 
         x"80", x"04", x"1E", x"00", x"00", x"00", x"24", x"10", x"20", x"80", 
         x"04", x"80", x"00", x"00", x"00", x"FF", x"18", x"00", x"00", x"00", 
         x"00", x"00", x"00", x"80", x"03", x"00", x"00", x"00", x"00", x"00", 
         x"00", x"00", x"80", x"03", x"00", x"00", x"80", x"00", x"28", x"20", 
         x"00", x"00", x"00", x"04", x"FF", x"FF", x"28", x"80", x"03", x"1E", 
         x"26", x"00", x"80", x"24", x"00", x"00", x"22", x"00", x"00", x"00", 
         x"00", x"00", x"99", x"90", x"80", x"04", x"1E", x"04", x"00", x"00", 
         x"00", x"00", x"00", x"28", x"00", x"00", x"FF", x"20", x"80", x"00", 
         x"00", x"80", x"90", x"00", x"04", x"80", x"04", x"00", x"FF", x"00", 
         x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"00", 
         x"00", x"00", x"00", x"00", x"A8", x"00", x"A0", x"00", x"00", x"01", 
         x"00", x"03", x"1E", x"98", x"1E", x"80", x"04", x"80", x"00", x"A9", 
         x"00", x"90", x"20", x"80", x"05", x"1E", x"00", x"00", x"00", x"00", 
         x"20", x"00", x"FF", x"20", x"80", x"00", x"00", x"80", x"90", x"00", 
         x"80", x"04", x"00", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", 
         x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"10", x"00", 
         x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"F0", 
         x"00", x"00", x"80", x"A0", x"88", x"1B", x"00", x"10", x"05", x"1B", 
         x"00", x"00", x"28", x"01", x"20", x"00", x"00", x"00", x"00", x"00", 
         x"20", x"FF", x"20", x"00", x"00", x"01", x"00", x"28", x"28", x"01", 
         x"20", x"00", x"20", x"00", x"20", x"28", x"00", x"01", x"00", x"FF", 
         x"00", x"20", x"F0", x"F0", x"00", x"00", x"00", x"98", x"80", x"1B", 
         x"00", x"05", x"1B", x"00", x"01", x"00", x"00", x"00", x"00", x"FF", 
         x"00", x"00", x"FF", x"20", x"00", x"00", x"01", x"00", x"28", x"01", 
         x"20", x"00", x"00", x"20", x"FF", x"01", x"00", x"00", x"FF", x"00", 
         x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
         x"00", x"00", x"05", x"88", x"05", x"80", x"FF", x"00", x"00", x"00", 
         x"00", x"01", x"00", x"00", x"03", x"1E", x"00", x"03", x"1E", x"05", 
         x"20", x"80", x"00", x"00", x"00", x"02", x"00", x"00", x"00", x"00", 
         x"00", x"00", x"00", x"FF", x"00", x"00", x"00", x"02", x"00", x"00", 
         x"00", x"FF", x"00", x"00", x"00", x"00", x"FF", x"05", x"20", x"05", 
         x"00", x"00", x"05", x"20", x"05", x"00", x"FF", x"00", x"00", x"00", 
         x"00", x"00", x"01", x"00", x"00", x"00", x"1E", x"1E", x"00", x"00", 
         x"00", x"00", x"03", x"80", x"00", x"00", x"00", x"10", x"00", x"00", 
         x"00", x"00", x"00", x"00", x"00", x"03", x"80", x"06", x"00", x"03", 
         x"1E", x"00", x"00", x"1E", x"00", x"00", x"02", x"00", x"00", x"00", 
         x"00", x"20", x"00", x"00", x"FF", x"00", x"80", x"00", x"00", x"00", 
         x"00", x"00", x"04", x"00", x"06", x"00", x"04", x"80", x"06", x"00", 
         x"04", x"80", x"06", x"00", x"FF", x"00", x"00", x"20", x"28", x"05", 
         x"00", x"00", x"00", x"06", x"00", x"05", x"00", x"09", x"07", x"07", 
         x"07", x"07", x"07", x"07", x"07", x"07", x"07", x"07", x"07", x"07", 
         x"07", x"07", x"07", x"07", x"07", x"07", x"07", x"07", x"07", x"07", 
         x"07", x"07", x"07", x"07", x"07", x"07", x"07", x"07", x"07", x"07", 
         x"07", x"07", x"07", x"07", x"07", x"07", x"07", x"07", x"07", x"07", 
         x"07", x"07", x"07", x"07", x"07", x"07", x"07", x"07", x"07", x"07", 
         x"07", x"07", x"07", x"07", x"07", x"07", x"07", x"07", x"07", x"07", 
         x"09", x"09", x"07", x"07", x"07", x"09", x"07", x"07", x"07", x"09", 
         x"07", x"09", x"07", x"07", x"07", x"07", x"0A", x"07", x"07", x"07", 
         x"07", x"0A", x"07", x"0A", x"09", x"07", x"07", x"07", x"07", x"07", 
         x"07", x"07", x"07", x"07", x"07", x"07", x"07", x"07", x"07", x"07", 
         x"07", x"07", x"07", x"07", x"07", x"07", x"07", x"07", x"07", x"07", 
         x"07", x"07", x"07", x"07", x"07", x"07", x"07", x"07", x"07", x"07", 
         x"07", x"07", x"07", x"07", x"07", x"07", x"07", x"07", x"07", x"07", 
         x"07", x"07", x"07", x"07", x"07", x"07", x"07", x"07", x"07", x"07", 
         x"07", x"07", x"07", x"07", x"07", x"07", x"09", x"09", x"07", x"07", 
         x"07", x"09", x"07", x"07", x"07", x"09", x"07", x"09", x"07", x"07", 
         x"07", x"07", x"09", x"07", x"07", x"07", x"07", x"09", x"07", x"09", 
         x"54", x"45", x"52", x"25", x"77", x"00", x"20", x"69", x"6F", x"6F", 
         x"72", x"2E", x"00", x"61", x"2E", x"00", x"65", x"65", x"79", x"6E", 
         x"74", x"2E", x"00", x"6C", x"20", x"67", x"2E", x"00", x"52", x"6D", 
         x"00", x"61", x"4D", x"72", x"00", x"52", x"61", x"00", x"61", x"67", 
         x"52", x"2E", x"61", x"55", x"61", x"00", x"6C", x"69", x"64", x"20", 
         x"00", x"69", x"67", x"72", x"63", x"69", x"74", x"73", x"73", x"20", 
         x"00", x"61", x"67", x"61", x"63", x"65", x"20", x"00", x"75", x"6E", 
         x"65", x"65", x"61", x"62", x"6B", x"00", x"75", x"6E", x"77", x"65", 
         x"20", x"73", x"00", x"61", x"62", x"6B", x"20", x"6B", x"00", x"61", 
         x"73", x"20", x"65", x"20", x"69", x"6C", x"6C", x"20", x"6F", x"00", 
         x"61", x"69", x"6E", x"20", x"6F", x"73", x"61", x"20", x"61", x"72", 
         x"61", x"00", x"61", x"69", x"6F", x"65", x"2C", x"74", x"67", x"74", 
         x"6F", x"20", x"00", x"B0", x"00", x"00", x"00", x"1D", x"1D", x"1D", 
         x"1B", x"1B", x"1C", x"00", x"1C", x"01", x"00", x"00", x"1C", x"00", 
         x"1C", x"00", x"1C", x"00", x"1C", x"00", x"1C", x"00", x"1C", x"00", 
         x"1D", x"00", x"1D", x"00", x"1D", x"32", x"00", x"1B", x"00", x"00", 
         x"32", x"00", x"1B", x"00", x"1D", x"62", x"00", x"1C", x"00", x"00", 
         x"62", x"00", x"1C", x"00", x"00", x"44", x"00", x"1C", x"00", x"1D", 
         x"1D", x"44", x"00", x"1C", x"00", x"1D", x"1D", others => x"00"
      ),
      2 => (
         x"1C", x"9C", x"1D", x"BD", x"02", x"42", x"03", x"63", x"40", x"42", 
         x"43", x"20", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
         x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
         x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
         x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"1A", x"40", 
         x"00", x"02", x"03", x"43", x"42", x"E0", x"42", x"03", x"02", x"43", 
         x"E0", x"00", x"02", x"82", x"A5", x"03", x"43", x"45", x"E0", x"00", 
         x"02", x"04", x"03", x"43", x"82", x"42", x"E0", x"00", x"02", x"82", 
         x"03", x"43", x"03", x"43", x"E0", x"00", x"03", x"05", x"65", x"62", 
         x"00", x"42", x"02", x"04", x"81", x"00", x"E0", x"00", x"02", x"E0", 
         x"00", x"04", x"E0", x"00", x"02", x"42", x"E0", x"42", x"84", x"02", 
         x"44", x"E0", x"00", x"C0", x"00", x"82", x"C6", x"A2", x"84", x"C0", 
         x"A5", x"E0", x"00", x"C0", x"05", x"05", x"C6", x"85", x"C0", x"84", 
         x"E0", x"00", x"82", x"00", x"40", x"00", x"00", x"42", x"82", x"63", 
         x"00", x"60", x"42", x"E0", x"42", x"E0", x"00", x"82", x"84", x"A2", 
         x"40", x"A5", x"E0", x"00", x"82", x"00", x"40", x"A5", x"45", x"84", 
         x"00", x"00", x"45", x"00", x"82", x"00", x"40", x"84", x"E0", x"00", 
         x"E0", x"00", x"E0", x"00", x"83", x"00", x"62", x"42", x"42", x"40", 
         x"02", x"62", x"00", x"60", x"05", x"00", x"84", x"65", x"00", x"60", 
         x"00", x"84", x"83", x"00", x"62", x"42", x"42", x"40", x"00", x"86", 
         x"00", x"C5", x"A2", x"42", x"40", x"84", x"00", x"86", x"02", x"02", 
         x"E2", x"45", x"C5", x"A6", x"C6", x"C0", x"84", x"04", x"64", x"00", 
         x"E0", x"00", x"E0", x"02", x"00", x"00", x"03", x"A3", x"03", x"A3", 
         x"A0", x"A3", x"A8", x"06", x"07", x"C4", x"A5", x"E5", x"65", x"63", 
         x"68", x"06", x"E0", x"60", x"03", x"A3", x"03", x"A3", x"A0", x"A7", 
         x"03", x"06", x"00", x"0A", x"63", x"E9", x"06", x"6A", x"E7", x"C4", 
         x"65", x"A5", x"A8", x"A9", x"00", x"A5", x"63", x"E5", x"06", x"6A", 
         x"E7", x"E0", x"40", x"82", x"00", x"02", x"62", x"02", x"62", x"02", 
         x"62", x"E0", x"82", x"04", x"04", x"05", x"05", x"04", x"03", x"00", 
         x"07", x"00", x"08", x"C8", x"00", x"45", x"05", x"05", x"63", x"04", 
         x"60", x"05", x"86", x"C7", x"00", x"45", x"05", x"05", x"63", x"04", 
         x"60", x"05", x"E0", x"00", x"A0", x"00", x"A0", x"00", x"E0", x"00", 
         x"05", x"80", x"00", x"A4", x"40", x"05", x"00", x"86", x"42", x"02", 
         x"A4", x"60", x"02", x"E0", x"00", x"00", x"04", x"E0", x"00", x"82", 
         x"00", x"40", x"42", x"82", x"00", x"40", x"42", x"82", x"02", x"E0", 
         x"82", x"E0", x"82", x"84", x"E0", x"85", x"84", x"82", x"40", x"A5", 
         x"84", x"A2", x"40", x"00", x"85", x"E0", x"00", x"02", x"43", x"40", 
         x"42", x"43", x"00", x"80", x"E0", x"80", x"05", x"A2", x"A5", x"43", 
         x"04", x"63", x"43", x"42", x"45", x"00", x"82", x"84", x"40", x"42", 
         x"44", x"00", x"82", x"00", x"40", x"42", x"E0", x"80", x"E0", x"82", 
         x"82", x"00", x"42", x"42", x"43", x"60", x"82", x"E0", x"00", x"00", 
         x"00", x"82", x"86", x"02", x"02", x"85", x"83", x"07", x"02", x"E2", 
         x"06", x"05", x"84", x"43", x"C5", x"63", x"63", x"A4", x"02", x"04", 
         x"BD", x"44", x"A5", x"67", x"BF", x"83", x"45", x"E0", x"00", x"00", 
         x"00", x"80", x"BF", x"00", x"E0", x"BD", x"BD", x"BF", x"B0", x"82", 
         x"00", x"40", x"90", x"44", x"00", x"10", x"02", x"00", x"40", x"44", 
         x"BF", x"B0", x"E0", x"BD", x"BD", x"B1", x"BF", x"B4", x"B3", x"B2", 
         x"B0", x"82", x"00", x"40", x"A0", x"13", x"12", x"80", x"73", x"14", 
         x"00", x"52", x"43", x"03", x"43", x"03", x"43", x"00", x"00", x"44", 
         x"02", x"00", x"40", x"10", x"03", x"43", x"43", x"60", x"03", x"03", 
         x"43", x"43", x"60", x"03", x"03", x"43", x"00", x"02", x"00", x"42", 
         x"42", x"43", x"60", x"10", x"02", x"42", x"42", x"00", x"40", x"00", 
         x"43", x"03", x"43", x"00", x"00", x"04", x"02", x"00", x"40", x"10", 
         x"BF", x"B4", x"B3", x"B2", x"B1", x"B0", x"E0", x"BD", x"03", x"04", 
         x"64", x"10", x"64", x"80", x"00", x"02", x"62", x"02", x"62", x"00", 
         x"20", x"00", x"85", x"00", x"40", x"00", x"00", x"02", x"00", x"42", 
         x"42", x"43", x"60", x"10", x"02", x"62", x"42", x"00", x"40", x"00", 
         x"00", x"80", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"80", 
         x"82", x"03", x"42", x"43", x"00", x"82", x"62", x"02", x"62", x"00", 
         x"20", x"00", x"85", x"00", x"40", x"00", x"00", x"00", x"04", x"00", 
         x"00", x"02", x"00", x"82", x"02", x"00", x"82", x"02", x"00", x"82", 
         x"00", x"80", x"02", x"00", x"82", x"02", x"00", x"82", x"02", x"00", 
         x"82", x"02", x"00", x"82", x"00", x"04", x"00", x"00", x"02", x"00", 
         x"82", x"02", x"00", x"82", x"02", x"00", x"82", x"00", x"80", x"02", 
         x"00", x"82", x"02", x"00", x"82", x"02", x"00", x"82", x"02", x"00", 
         x"82", x"00", x"20", x"00", x"00", x"00", x"04", x"00", x"00", x"00", 
         x"24", x"00", x"00", x"02", x"43", x"82", x"03", x"84", x"E0", x"83", 
         x"BD", x"B5", x"15", x"B4", x"B3", x"B2", x"B1", x"BF", x"B0", x"00", 
         x"B5", x"12", x"13", x"14", x"42", x"23", x"50", x"02", x"00", x"82", 
         x"13", x"90", x"60", x"00", x"14", x"00", x"20", x"00", x"00", x"00", 
         x"82", x"83", x"02", x"02", x"A4", x"02", x"82", x"43", x"02", x"B1", 
         x"52", x"40", x"60", x"42", x"31", x"50", x"02", x"23", x"00", x"82", 
         x"13", x"90", x"B1", x"20", x"BF", x"A0", x"B4", x"B5", x"B3", x"B2", 
         x"B1", x"B0", x"E0", x"BD", x"00", x"00", x"B1", x"50", x"00", x"31", 
         x"BD", x"B1", x"B1", x"B2", x"BF", x"B0", x"20", x"92", x"00", x"40", 
         x"00", x"10", x"02", x"51", x"40", x"40", x"BF", x"B2", x"B1", x"B0", 
         x"E0", x"BD", x"BD", x"B3", x"B1", x"BF", x"B7", x"B6", x"B5", x"B4", 
         x"B2", x"B0", x"83", x"B4", x"A2", x"83", x"97", x"A3", x"94", x"80", 
         x"A0", x"95", x"94", x"60", x"E2", x"A2", x"B5", x"F6", x"B5", x"00", 
         x"00", x"F7", x"00", x"A2", x"44", x"00", x"10", x"A2", x"04", x"C2", 
         x"00", x"45", x"22", x"10", x"02", x"40", x"00", x"90", x"A5", x"00", 
         x"A0", x"02", x"02", x"22", x"52", x"00", x"44", x"00", x"00", x"23", 
         x"00", x"70", x"04", x"65", x"64", x"00", x"A2", x"00", x"04", x"44", 
         x"00", x"10", x"A2", x"04", x"E2", x"00", x"45", x"00", x"04", x"64", 
         x"65", x"00", x"10", x"22", x"00", x"02", x"40", x"90", x"BF", x"B7", 
         x"B6", x"B5", x"B4", x"B3", x"B2", x"B1", x"B0", x"E0", x"BD", x"BD", 
         x"B0", x"84", x"F0", x"BF", x"B2", x"B1", x"B2", x"00", x"D1", x"05", 
         x"40", x"00", x"A5", x"20", x"BF", x"B2", x"B1", x"B0", x"00", x"BD", 
         x"BD", x"BF", x"B4", x"B0", x"B3", x"80", x"B2", x"B1", x"82", x"91", 
         x"05", x"84", x"13", x"12", x"00", x"22", x"04", x"05", x"00", x"31", 
         x"07", x"06", x"04", x"00", x"05", x"05", x"04", x"A5", x"00", x"A5", 
         x"07", x"06", x"04", x"00", x"05", x"04", x"05", x"84", x"A5", x"A5", 
         x"00", x"84", x"04", x"00", x"31", x"05", x"04", x"A5", x"00", x"A5", 
         x"07", x"04", x"05", x"00", x"06", x"14", x"00", x"94", x"94", x"91", 
         x"40", x"72", x"52", x"52", x"04", x"00", x"80", x"00", x"04", x"80", 
         x"40", x"00", x"94", x"94", x"00", x"04", x"91", x"40", x"00", x"04", 
         x"00", x"20", x"07", x"05", x"06", x"00", x"04", x"00", x"00", x"BF", 
         x"B4", x"B3", x"B2", x"B1", x"B0", x"04", x"00", x"00", x"BD", x"BD", 
         x"B0", x"80", x"84", x"BF", x"00", x"B1", x"42", x"00", x"51", x"05", 
         x"B1", x"03", x"62", x"05", x"51", x"85", x"05", x"50", x"BF", x"B1", 
         x"B0", x"40", x"BD", x"00", x"65", x"BD", x"B1", x"80", x"A4", x"B0", 
         x"BF", x"00", x"A0", x"03", x"26", x"24", x"05", x"64", x"C5", x"31", 
         x"84", x"A5", x"22", x"A5", x"84", x"00", x"23", x"00", x"04", x"04", 
         x"00", x"00", x"25", x"BF", x"B1", x"B0", x"04", x"A5", x"00", x"BD", 
         x"BD", x"BF", x"B0", x"A0", x"02", x"A3", x"86", x"85", x"C3", x"A2", 
         x"84", x"A5", x"84", x"00", x"A5", x"05", x"00", x"04", x"02", x"05", 
         x"A2", x"BF", x"B0", x"04", x"A5", x"00", x"BD", x"BD", x"B1", x"BF", 
         x"B3", x"B2", x"B0", x"86", x"00", x"C0", x"80", x"00", x"12", x"00", 
         x"13", x"00", x"00", x"26", x"10", x"10", x"06", x"40", x"00", x"02", 
         x"02", x"22", x"42", x"20", x"43", x"00", x"72", x"40", x"60", x"00", 
         x"73", x"00", x"00", x"20", x"10", x"26", x"10", x"06", x"40", x"02", 
         x"BF", x"B3", x"B2", x"B1", x"B0", x"E0", x"BD", x"00", x"10", x"26", 
         x"00", x"10", x"A3", x"A2", x"63", x"43", x"42", x"00", x"A2", x"00", 
         x"A0", x"A2", x"00", x"40", x"42", x"00", x"A2", x"A2", x"00", x"42", 
         x"00", x"A2", x"BD", x"BF", x"00", x"00", x"43", x"60", x"42", x"40", 
         x"84", x"BF", x"00", x"E0", x"BD", x"BF", x"00", x"BD", x"BF", x"84", 
         x"00", x"BD", x"BD", x"B4", x"14", x"BF", x"B0", x"B3", x"B2", x"00", 
         x"B1", x"00", x"84", x"84", x"00", x"85", x"84", x"85", x"80", x"00", 
         x"10", x"00", x"10", x"11", x"10", x"00", x"51", x"02", x"42", x"22", 
         x"40", x"84", x"00", x"85", x"11", x"84", x"85", x"80", x"00", x"73", 
         x"00", x"00", x"92", x"60", x"00", x"00", x"10", x"10", x"40", x"85", 
         x"00", x"82", x"00", x"10", x"42", x"40", x"13", x"BF", x"B4", x"B3", 
         x"B2", x"B1", x"B0", x"84", x"00", x"BD", x"BF", x"B4", x"B3", x"B2", 
         x"B1", x"B0", x"84", x"00", x"BD", x"12", x"00", x"13", x"51", x"00", 
         x"A5", x"00", x"10", x"00", x"52", x"13", x"51", x"85", x"00", x"84", 
         x"11", x"00", x"80", x"11", x"00", x"84", x"11", x"00", x"84", x"00", 
         x"24", x"20", x"11", x"60", x"00", x"00", x"94", x"00", x"10", x"11", 
         x"00", x"00", x"00", x"40", x"00", x"04", x"12", x"80", x"82", x"00", 
         x"42", x"85", x"13", x"10", x"00", x"82", x"00", x"00", x"11", x"00", 
         x"BF", x"B4", x"B3", x"B2", x"B1", x"B0", x"00", x"BD", x"BD", x"B0", 
         x"10", x"BF", x"B5", x"B4", x"A0", x"B3", x"80", x"B6", x"B2", x"00", 
         x"B1", x"00", x"04", x"15", x"04", x"85", x"00", x"80", x"60", x"15", 
         x"16", x"A0", x"11", x"00", x"00", x"D6", x"10", x"13", x"31", x"00", 
         x"14", x"22", x"12", x"C0", x"82", x"00", x"42", x"85", x"15", x"10", 
         x"82", x"00", x"31", x"13", x"00", x"BF", x"B6", x"B5", x"B4", x"B3", 
         x"B2", x"B1", x"B0", x"E0", x"BD", x"BD", x"B2", x"92", x"92", x"BE", 
         x"BF", x"B7", x"B6", x"B5", x"B4", x"B3", x"B1", x"B0", x"40", x"80", 
         x"02", x"16", x"80", x"00", x"00", x"53", x"15", x"17", x"00", x"D6", 
         x"00", x"00", x"40", x"00", x"60", x"35", x"22", x"51", x"10", x"12", 
         x"02", x"20", x"00", x"85", x"04", x"00", x"A5", x"10", x"B7", x"00", 
         x"C0", x"00", x"00", x"94", x"60", x"40", x"10", x"00", x"94", x"12", 
         x"11", x"02", x"1E", x"C2", x"15", x"02", x"11", x"00", x"00", x"52", 
         x"14", x"00", x"B5", x"C5", x"00", x"00", x"14", x"02", x"50", x"31", 
         x"20", x"DE", x"00", x"40", x"65", x"04", x"00", x"A5", x"C0", x"00", 
         x"A0", x"C5", x"73", x"40", x"31", x"00", x"73", x"10", x"20", x"DE", 
         x"BF", x"BE", x"B7", x"B6", x"B5", x"B4", x"B3", x"B2", x"B1", x"B0", 
         x"E0", x"BD", x"00", x"00", x"00", x"00", x"BD", x"BF", x"B3", x"B2", 
         x"B1", x"00", x"B0", x"04", x"00", x"84", x"04", x"00", x"84", x"00", 
         x"00", x"00", x"11", x"12", x"13", x"00", x"00", x"42", x"00", x"51", 
         x"00", x"52", x"00", x"53", x"00", x"00", x"00", x"00", x"00", x"42", 
         x"00", x"51", x"00", x"02", x"40", x"00", x"10", x"00", x"00", x"00", 
         x"00", x"10", x"00", x"00", x"00", x"00", x"BD", x"BF", x"B4", x"B3", 
         x"B2", x"B1", x"00", x"B0", x"00", x"00", x"02", x"03", x"61", x"42", 
         x"40", x"11", x"00", x"84", x"00", x"00", x"BF", x"00", x"B4", x"B3", 
         x"B2", x"B1", x"B0", x"E0", x"BD", x"00", x"84", x"00", x"00", x"00", 
         x"24", x"10", x"12", x"31", x"14", x"13", x"00", x"00", x"42", x"00", 
         x"50", x"20", x"52", x"00", x"54", x"00", x"82", x"00", x"53", x"00", 
         x"40", x"03", x"00", x"00", x"00", x"00", x"00", x"85", x"00", x"00", 
         x"00", x"85", x"00", x"00", x"43", x"00", x"00", x"00", x"40", x"00", 
         x"04", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
         x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
         x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
         x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
         x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
         x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
         x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
         x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
         x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
         x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
         x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
         x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
         x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
         x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
         x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
         x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
         x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
         x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
         x"41", x"20", x"4F", x"79", x"24", x"00", x"78", x"6F", x"42", x"6C", 
         x"65", x"30", x"32", x"74", x"20", x"00", x"69", x"6D", x"72", x"6F", 
         x"6E", x"2E", x"00", x"70", x"64", x"61", x"2E", x"00", x"44", x"65", 
         x"79", x"6C", x"20", x"6F", x"00", x"44", x"6F", x"00", x"6F", x"6E", 
         x"44", x"2E", x"6D", x"20", x"6F", x"00", x"70", x"64", x"20", x"61", 
         x"2E", x"61", x"6E", x"6F", x"6E", x"6D", x"20", x"6E", x"73", x"6E", 
         x"2E", x"72", x"6E", x"6C", x"20", x"74", x"73", x"2E", x"6F", x"20", 
         x"20", x"73", x"6C", x"20", x"63", x"00", x"6F", x"20", x"20", x"74", 
         x"6F", x"61", x"00", x"6C", x"20", x"63", x"73", x"63", x"2E", x"6D", 
         x"20", x"65", x"63", x"73", x"61", x"62", x"66", x"68", x"6D", x"2E", 
         x"6C", x"20", x"69", x"6E", x"72", x"75", x"74", x"2E", x"65", x"20", 
         x"74", x"2E", x"6C", x"20", x"6E", x"72", x"79", x"6C", x"75", x"69", 
         x"68", x"64", x"2E", x"B9", x"00", x"00", x"00", x"00", x"00", x"00", 
         x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
         x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
         x"00", x"00", x"00", x"00", x"00", x"0C", x"00", x"00", x"00", x"00", 
         x"0C", x"00", x"00", x"00", x"00", x"11", x"00", x"00", x"00", x"00", 
         x"01", x"00", x"00", x"00", x"00", x"0C", x"00", x"00", x"00", x"00", 
         x"00", x"0C", x"00", x"00", x"00", x"00", x"00", others => x"00"
      ),
      3 => (
         x"3C", x"27", x"3C", x"27", x"3C", x"24", x"3C", x"24", x"AC", x"24", 
         x"00", x"14", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
         x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
         x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
         x"00", x"00", x"0C", x"00", x"00", x"08", x"00", x"00", x"3C", x"03", 
         x"00", x"3C", x"24", x"A0", x"90", x"03", x"30", x"24", x"3C", x"A0", 
         x"03", x"00", x"3C", x"00", x"30", x"24", x"A0", x"A0", x"03", x"00", 
         x"3C", x"00", x"24", x"A0", x"00", x"8C", x"03", x"00", x"3C", x"00", 
         x"24", x"A0", x"24", x"A0", x"03", x"00", x"3C", x"24", x"A0", x"90", 
         x"00", x"30", x"00", x"00", x"04", x"00", x"03", x"00", x"8C", x"03", 
         x"00", x"AC", x"03", x"00", x"3C", x"8C", x"03", x"30", x"30", x"3C", 
         x"AC", x"03", x"00", x"10", x"00", x"80", x"24", x"A0", x"24", x"14", 
         x"24", x"03", x"00", x"10", x"00", x"00", x"24", x"A0", x"14", x"24", 
         x"03", x"00", x"90", x"00", x"10", x"00", x"00", x"24", x"00", x"90", 
         x"00", x"14", x"24", x"03", x"24", x"03", x"00", x"90", x"24", x"A0", 
         x"14", x"24", x"03", x"00", x"90", x"00", x"10", x"30", x"10", x"24", 
         x"08", x"00", x"10", x"00", x"90", x"00", x"14", x"24", x"03", x"00", 
         x"03", x"00", x"03", x"00", x"90", x"00", x"24", x"30", x"2C", x"14", 
         x"24", x"10", x"00", x"10", x"24", x"08", x"24", x"10", x"00", x"10", 
         x"00", x"24", x"90", x"00", x"24", x"30", x"2C", x"10", x"00", x"90", 
         x"00", x"24", x"30", x"2C", x"10", x"24", x"00", x"90", x"00", x"00", 
         x"00", x"00", x"24", x"30", x"2C", x"14", x"24", x"24", x"10", x"00", 
         x"03", x"00", x"03", x"00", x"08", x"00", x"24", x"A0", x"24", x"A0", 
         x"00", x"24", x"24", x"3C", x"24", x"00", x"2C", x"00", x"A0", x"24", 
         x"14", x"00", x"03", x"A0", x"24", x"A0", x"24", x"A0", x"00", x"24", 
         x"24", x"3C", x"08", x"24", x"24", x"A0", x"00", x"10", x"24", x"00", 
         x"00", x"30", x"2C", x"24", x"15", x"24", x"24", x"A0", x"00", x"14", 
         x"24", x"03", x"A0", x"8F", x"00", x"00", x"00", x"00", x"00", x"00", 
         x"00", x"03", x"AF", x"00", x"00", x"00", x"00", x"00", x"24", x"00", 
         x"24", x"08", x"24", x"14", x"00", x"00", x"00", x"00", x"24", x"00", 
         x"10", x"00", x"30", x"14", x"00", x"00", x"00", x"00", x"24", x"00", 
         x"14", x"00", x"03", x"00", x"04", x"00", x"14", x"00", x"03", x"00", 
         x"00", x"04", x"00", x"00", x"10", x"00", x"00", x"00", x"24", x"00", 
         x"00", x"14", x"00", x"03", x"00", x"08", x"00", x"03", x"00", x"93", 
         x"00", x"14", x"24", x"93", x"00", x"10", x"24", x"A3", x"24", x"03", 
         x"A3", x"03", x"A3", x"A3", x"03", x"A3", x"30", x"2C", x"10", x"30", 
         x"A3", x"2C", x"10", x"00", x"A3", x"03", x"00", x"3C", x"24", x"A4", 
         x"24", x"14", x"00", x"A3", x"03", x"A3", x"3C", x"24", x"24", x"94", 
         x"3C", x"30", x"A4", x"24", x"14", x"00", x"24", x"24", x"A4", x"24", 
         x"14", x"00", x"93", x"00", x"14", x"24", x"03", x"A3", x"03", x"A3", 
         x"93", x"00", x"24", x"30", x"2C", x"10", x"A3", x"03", x"00", x"08", 
         x"00", x"93", x"93", x"00", x"00", x"93", x"93", x"01", x"00", x"00", 
         x"00", x"00", x"30", x"00", x"00", x"24", x"30", x"00", x"00", x"3C", 
         x"27", x"00", x"30", x"2C", x"AF", x"A3", x"A4", x"14", x"00", x"0C", 
         x"00", x"A3", x"8F", x"00", x"03", x"27", x"27", x"AF", x"AF", x"80", 
         x"00", x"10", x"24", x"30", x"0C", x"26", x"82", x"00", x"14", x"30", 
         x"8F", x"8F", x"03", x"27", x"27", x"AF", x"AF", x"AF", x"AF", x"AF", 
         x"AF", x"80", x"00", x"10", x"00", x"3C", x"3C", x"00", x"26", x"3C", 
         x"08", x"26", x"10", x"24", x"10", x"24", x"10", x"00", x"0C", x"30", 
         x"82", x"00", x"10", x"26", x"24", x"10", x"28", x"14", x"24", x"24", 
         x"10", x"28", x"10", x"24", x"24", x"14", x"00", x"92", x"00", x"24", 
         x"30", x"2C", x"10", x"26", x"00", x"02", x"8C", x"00", x"00", x"00", 
         x"10", x"24", x"14", x"00", x"0C", x"24", x"82", x"00", x"14", x"26", 
         x"8F", x"8F", x"8F", x"8F", x"8F", x"8F", x"03", x"27", x"82", x"24", 
         x"10", x"26", x"28", x"14", x"00", x"24", x"10", x"24", x"14", x"00", 
         x"02", x"0C", x"26", x"0C", x"00", x"08", x"00", x"92", x"00", x"24", 
         x"30", x"2C", x"10", x"26", x"00", x"02", x"8C", x"00", x"00", x"00", 
         x"08", x"A3", x"0C", x"00", x"08", x"00", x"0C", x"00", x"08", x"A3", 
         x"93", x"24", x"24", x"00", x"08", x"A3", x"10", x"24", x"14", x"00", 
         x"02", x"0C", x"26", x"0C", x"00", x"08", x"00", x"0C", x"24", x"08", 
         x"00", x"24", x"08", x"A3", x"24", x"08", x"A3", x"24", x"08", x"A3", 
         x"08", x"A3", x"24", x"08", x"A3", x"24", x"08", x"A3", x"24", x"08", 
         x"A3", x"24", x"08", x"A3", x"0C", x"24", x"08", x"00", x"24", x"08", 
         x"A3", x"24", x"08", x"A3", x"24", x"08", x"A3", x"08", x"A3", x"24", 
         x"08", x"A3", x"24", x"08", x"A3", x"24", x"08", x"A3", x"24", x"08", 
         x"A3", x"0C", x"02", x"08", x"00", x"0C", x"24", x"08", x"00", x"0C", 
         x"32", x"08", x"00", x"3C", x"8C", x"27", x"00", x"A3", x"03", x"A3", 
         x"27", x"AF", x"3C", x"AF", x"AF", x"AF", x"AF", x"AF", x"AF", x"00", 
         x"26", x"3C", x"24", x"24", x"8E", x"2A", x"30", x"00", x"02", x"A3", 
         x"12", x"A3", x"10", x"00", x"16", x"00", x"12", x"00", x"0C", x"00", 
         x"93", x"93", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"02", 
         x"00", x"A4", x"A0", x"8E", x"26", x"30", x"00", x"2A", x"02", x"A3", 
         x"16", x"A3", x"02", x"A2", x"8F", x"02", x"8F", x"8F", x"8F", x"8F", 
         x"8F", x"8F", x"03", x"27", x"0C", x"00", x"02", x"A0", x"08", x"26", 
         x"27", x"AF", x"30", x"AF", x"AF", x"AF", x"12", x"30", x"00", x"02", 
         x"0C", x"26", x"32", x"00", x"14", x"02", x"8F", x"8F", x"8F", x"8F", 
         x"03", x"27", x"27", x"AF", x"AF", x"AF", x"AF", x"AF", x"AF", x"AF", 
         x"AF", x"AF", x"90", x"90", x"90", x"02", x"90", x"90", x"26", x"00", 
         x"00", x"90", x"32", x"10", x"02", x"02", x"26", x"26", x"32", x"00", 
         x"08", x"26", x"0C", x"AF", x"8E", x"0C", x"26", x"8F", x"24", x"02", 
         x"0C", x"30", x"92", x"32", x"02", x"10", x"00", x"02", x"30", x"0C", 
         x"02", x"26", x"00", x"02", x"8C", x"00", x"8E", x"0C", x"00", x"92", 
         x"00", x"14", x"24", x"92", x"92", x"0C", x"AF", x"0C", x"24", x"8E", 
         x"0C", x"26", x"8F", x"24", x"02", x"0C", x"30", x"0C", x"24", x"92", 
         x"92", x"0C", x"32", x"92", x"00", x"02", x"14", x"02", x"8F", x"8F", 
         x"8F", x"8F", x"8F", x"8F", x"8F", x"8F", x"8F", x"03", x"27", x"27", 
         x"AF", x"30", x"30", x"AF", x"AF", x"AF", x"30", x"0C", x"30", x"26", 
         x"02", x"0C", x"30", x"02", x"8F", x"8F", x"8F", x"8F", x"08", x"27", 
         x"27", x"AF", x"AF", x"AF", x"AF", x"00", x"AF", x"AF", x"90", x"90", 
         x"92", x"90", x"92", x"92", x"0C", x"02", x"92", x"92", x"0C", x"26", 
         x"92", x"24", x"24", x"0C", x"24", x"92", x"92", x"24", x"0C", x"30", 
         x"92", x"24", x"24", x"0C", x"24", x"92", x"92", x"24", x"24", x"30", 
         x"0C", x"30", x"8E", x"0C", x"32", x"92", x"92", x"24", x"0C", x"30", 
         x"92", x"24", x"24", x"0C", x"24", x"92", x"00", x"26", x"32", x"02", 
         x"10", x"02", x"26", x"32", x"92", x"0C", x"02", x"0C", x"24", x"02", 
         x"02", x"0C", x"26", x"32", x"0C", x"24", x"02", x"14", x"00", x"92", 
         x"0C", x"02", x"92", x"24", x"24", x"0C", x"24", x"0C", x"02", x"8F", 
         x"8F", x"8F", x"8F", x"8F", x"8F", x"24", x"00", x"08", x"27", x"27", 
         x"AF", x"00", x"8C", x"AF", x"0C", x"AF", x"24", x"0C", x"30", x"24", 
         x"00", x"3C", x"24", x"00", x"A0", x"00", x"00", x"AC", x"8F", x"8F", 
         x"8F", x"00", x"27", x"08", x"A0", x"27", x"AF", x"00", x"8C", x"AF", 
         x"AF", x"0C", x"00", x"92", x"92", x"92", x"92", x"00", x"00", x"92", 
         x"24", x"24", x"02", x"30", x"30", x"0C", x"02", x"0C", x"24", x"8E", 
         x"0C", x"00", x"26", x"8F", x"8F", x"8F", x"24", x"30", x"08", x"27", 
         x"27", x"AF", x"AF", x"00", x"92", x"90", x"90", x"90", x"00", x"00", 
         x"24", x"24", x"30", x"0C", x"30", x"92", x"0C", x"24", x"8E", x"24", 
         x"00", x"8F", x"8F", x"24", x"30", x"08", x"27", x"27", x"AF", x"AF", 
         x"AF", x"AF", x"AF", x"90", x"00", x"10", x"00", x"00", x"24", x"08", 
         x"24", x"0C", x"00", x"92", x"26", x"32", x"02", x"10", x"00", x"26", 
         x"00", x"02", x"8C", x"02", x"90", x"00", x"10", x"00", x"10", x"00", 
         x"14", x"00", x"0C", x"02", x"26", x"92", x"32", x"02", x"14", x"26", 
         x"8F", x"8F", x"8F", x"8F", x"8F", x"03", x"27", x"0C", x"26", x"92", 
         x"08", x"32", x"90", x"90", x"24", x"10", x"24", x"08", x"A0", x"08", 
         x"A0", x"90", x"00", x"10", x"24", x"08", x"A0", x"90", x"00", x"24", 
         x"08", x"A0", x"27", x"AF", x"0C", x"00", x"30", x"14", x"30", x"14", 
         x"27", x"8F", x"00", x"03", x"27", x"8F", x"08", x"27", x"8F", x"27", 
         x"08", x"27", x"27", x"AF", x"3C", x"AF", x"AF", x"AF", x"AF", x"0C", 
         x"AF", x"0C", x"26", x"26", x"0C", x"27", x"26", x"27", x"AF", x"0C", 
         x"24", x"0C", x"26", x"00", x"32", x"16", x"00", x"3C", x"24", x"02", 
         x"10", x"26", x"0C", x"27", x"00", x"26", x"27", x"AF", x"0C", x"26", 
         x"00", x"08", x"26", x"10", x"00", x"0C", x"00", x"00", x"02", x"27", 
         x"0C", x"AF", x"0C", x"26", x"30", x"10", x"02", x"8F", x"8F", x"8F", 
         x"8F", x"8F", x"8F", x"27", x"08", x"27", x"8F", x"8F", x"8F", x"8F", 
         x"8F", x"8F", x"27", x"08", x"27", x"24", x"00", x"24", x"02", x"02", 
         x"30", x"0C", x"26", x"0C", x"26", x"16", x"02", x"27", x"0C", x"26", 
         x"00", x"0C", x"AF", x"00", x"0C", x"30", x"00", x"0C", x"30", x"0C", 
         x"32", x"12", x"00", x"02", x"00", x"08", x"26", x"0C", x"26", x"12", 
         x"00", x"0C", x"00", x"00", x"0C", x"26", x"16", x"02", x"8F", x"00", 
         x"24", x"27", x"02", x"26", x"0C", x"AF", x"0C", x"00", x"16", x"00", 
         x"8F", x"8F", x"8F", x"8F", x"8F", x"8F", x"08", x"27", x"27", x"AF", 
         x"3C", x"AF", x"AF", x"AF", x"00", x"AF", x"00", x"AF", x"AF", x"0C", 
         x"AF", x"0C", x"26", x"00", x"26", x"27", x"0C", x"AF", x"12", x"00", 
         x"3C", x"02", x"3C", x"00", x"08", x"26", x"26", x"12", x"26", x"0C", 
         x"02", x"AE", x"16", x"02", x"8F", x"00", x"24", x"27", x"02", x"26", 
         x"AF", x"0C", x"26", x"16", x"00", x"8F", x"8F", x"8F", x"8F", x"8F", 
         x"8F", x"8F", x"8F", x"03", x"27", x"27", x"AF", x"24", x"00", x"AF", 
         x"AF", x"AF", x"AF", x"AF", x"AF", x"AF", x"AF", x"AF", x"10", x"00", 
         x"3C", x"3C", x"00", x"00", x"00", x"24", x"24", x"3C", x"08", x"26", 
         x"0C", x"00", x"00", x"0C", x"02", x"12", x"26", x"30", x"26", x"12", 
         x"3C", x"16", x"02", x"26", x"24", x"0C", x"30", x"00", x"00", x"0C", 
         x"02", x"0C", x"02", x"26", x"02", x"00", x"26", x"0C", x"32", x"16", 
         x"24", x"3C", x"00", x"03", x"3C", x"3C", x"24", x"00", x"00", x"24", 
         x"24", x"08", x"26", x"8F", x"0C", x"00", x"12", x"26", x"30", x"26", 
         x"12", x"27", x"16", x"02", x"26", x"24", x"0C", x"30", x"03", x"0C", 
         x"02", x"8F", x"26", x"02", x"26", x"0C", x"32", x"24", x"16", x"27", 
         x"8F", x"8F", x"8F", x"8F", x"8F", x"8F", x"8F", x"8F", x"8F", x"8F", 
         x"03", x"27", x"08", x"00", x"08", x"00", x"27", x"AF", x"AF", x"AF", 
         x"AF", x"0C", x"AF", x"3C", x"0C", x"24", x"3C", x"0C", x"24", x"0C", 
         x"00", x"00", x"24", x"24", x"24", x"0C", x"00", x"90", x"00", x"10", 
         x"00", x"10", x"00", x"14", x"00", x"0C", x"00", x"0C", x"00", x"90", 
         x"00", x"14", x"00", x"2E", x"14", x"00", x"26", x"0C", x"02", x"08", 
         x"00", x"26", x"0C", x"02", x"08", x"00", x"27", x"AF", x"AF", x"AF", 
         x"AF", x"AF", x"0C", x"AF", x"0C", x"00", x"00", x"00", x"04", x"30", 
         x"10", x"3C", x"0C", x"27", x"0C", x"00", x"8F", x"00", x"8F", x"8F", 
         x"8F", x"8F", x"8F", x"03", x"27", x"0C", x"27", x"08", x"00", x"0C", 
         x"26", x"24", x"24", x"26", x"24", x"24", x"0C", x"00", x"90", x"00", 
         x"10", x"02", x"10", x"00", x"14", x"00", x"93", x"00", x"10", x"00", 
         x"14", x"24", x"0C", x"00", x"08", x"00", x"0C", x"27", x"08", x"00", 
         x"0C", x"27", x"08", x"00", x"14", x"00", x"0C", x"00", x"00", x"0C", 
         x"24", x"0C", x"00", x"08", x"00", x"0C", x"00", x"00", x"00", x"00", 
         x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
         x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
         x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
         x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
         x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
         x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
         x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
         x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
         x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
         x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
         x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
         x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
         x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
         x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
         x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
         x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
         x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
         x"46", x"4C", x"52", x"24", x"3A", x"00", x"25", x"76", x"20", x"74", 
         x"64", x"76", x"2E", x"53", x"74", x"2E", x"56", x"20", x"6F", x"63", 
         x"65", x"20", x"00", x"55", x"61", x"6D", x"20", x"00", x"44", x"4D", 
         x"72", x"46", x"68", x"6D", x"00", x"44", x"4C", x"00", x"4C", x"69", 
         x"44", x"2E", x"49", x"65", x"6C", x"00", x"55", x"61", x"67", x"74", 
         x"2E", x"57", x"69", x"66", x"69", x"6D", x"67", x"61", x"69", x"6F", 
         x"2E", x"45", x"69", x"66", x"68", x"6E", x"74", x"2E", x"43", x"64", 
         x"74", x"61", x"66", x"68", x"6F", x"00", x"43", x"64", x"74", x"69", 
         x"74", x"6C", x"2E", x"46", x"68", x"6F", x"69", x"6F", x"64", x"49", 
         x"65", x"7A", x"78", x"64", x"76", x"61", x"20", x"73", x"65", x"79", 
         x"46", x"68", x"20", x"61", x"72", x"6F", x"73", x"65", x"6C", x"65", 
         x"73", x"74", x"46", x"68", x"20", x"20", x"64", x"61", x"6F", x"20", 
         x"73", x"6C", x"65", x"12", x"07", x"01", x"03", x"00", x"00", x"00", 
         x"00", x"00", x"00", x"00", x"00", x"02", x"00", x"00", x"00", x"00", 
         x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
         x"00", x"00", x"00", x"00", x"00", x"19", x"04", x"00", x"01", x"00", 
         x"19", x"07", x"00", x"01", x"00", x"01", x"06", x"00", x"00", x"00", 
         x"01", x"06", x"00", x"00", x"00", x"10", x"07", x"00", x"02", x"00", 
         x"00", x"10", x"07", x"00", x"02", x"00", x"00", others => x"00"
      )
   );

end data;